
module tb_ROC_RV32_program;
	timeunit 1ns;
	timeprecision 1ps;

	logic clk;
	logic rst_n;

	soc #(
		.ADDR_WIDTH_I(10),
		.DATA_WIDTH_I(32),
		.ADDR_WIDTH_D(10),
		.DATA_WIDTH_D(32)
	) dut (
		.clk(clk),
		.rst_n(rst_n),
		.imem_b_en(1'b0),
		.imem_b_we(1'b0),
		.imem_b_wstrb(4'b0000),
		.imem_b_addr('0),
		.imem_b_wdata('0),
		.imem_b_rdata(),
		.dmem_b_en(1'b0),
		.dmem_b_we(1'b0),
		.dmem_b_wstrb(4'b0000),
		.dmem_b_addr('0),
		.dmem_b_wdata('0),
		.dmem_b_rdata()
	);

	initial clk = 1'b0;
	always #5 clk = ~clk;

	task automatic reset_dut();
		rst_n = 1'b0;
		repeat (5) @(posedge clk);
		rst_n = 1'b1;
		repeat (2) @(posedge clk);
	endtask

	int unsigned cycles;
	int unsigned store_count;
	logic        saw_store_to_word0;
	logic        saw_fail_signature;
	logic [31:0] last_word0_wdata;
	int unsigned stop_addr_word;
	int unsigned max_cycles;
	logic [31:0] stop_wdata;
	bit          use_stop_wdata;
	string imem_path;
	integer fd;

	task automatic dump_dmem();
		$display("---- DMEM DUMP (word-addressed) ----");
		for (int i = 0; i < 100; i++) begin
			$display("dmem[%0d]=0x%08x", i, dut.data_memory.data_memory.mem[i]);
		end
		$display("----------------------------------");
	endtask

	initial begin
		rst_n = 1'b0;

		// Stop condition configuration:
		// - default: stop on an exact store of 0xDEADBEEF to dmem[word 0]
		// - optional: stop on an exact store value with +STOP_WDATA=<hex>
		// - optional: change stop address with +STOP_ADDR=<decimal word index>
		// - optional: change timeout with +MAX_CYCLES=<decimal>
		stop_addr_word = 0;
		max_cycles = 5_000_000;
		stop_wdata = 32'hDEAD_BEEF;
		use_stop_wdata = 1'b1;
		void'($value$plusargs("STOP_ADDR=%d", stop_addr_word));
		void'($value$plusargs("MAX_CYCLES=%d", max_cycles));
		if ($value$plusargs("STOP_WDATA=%h", stop_wdata)) begin
			use_stop_wdata = 1'b1;
		end

		// Clear dmem
		for (int i = 0; i < 18; i++) begin
			dut.data_memory.data_memory.mem[i] = 32'h0000_0000;
		end

		// Load program into imem (generated by `make`).
		// Note: Questa runs from ./questasim (see run_sim.tcl), so we try paths relative to that.
		imem_path = "sw/imem.dat";
		fd = $fopen(imem_path, "r");
		if (fd == 0) begin
			imem_path = "../sw/imem.dat";
			fd = $fopen(imem_path, "r");
		end
		if (fd == 0) begin
			$fatal(1, "Failed to open sw/imem.dat (tried sw/imem.dat and ../sw/imem.dat)");
		end
		$fclose(fd);
		$display("[TB] Loading IMEM from: %s", imem_path);
		$readmemh(imem_path, dut.instruction_memory.data_memory.mem);

		reset_dut();

		cycles = 0;
		store_count = 0;
		saw_store_to_word0 = 1'b0;
		saw_fail_signature = 1'b0;
		last_word0_wdata = 32'h0000_0000;

		// Stop when the program signals completion by writing the signature.
		// Override with +STOP_WDATA=... and/or +STOP_ADDR=... if needed.
		while (!saw_store_to_word0 && cycles < max_cycles) begin
			@(posedge clk);
			cycles++;

			if (rst_n && dut.cpu_core.cpu_state == 3'd4) begin
				$display("[WB] pc=0x%08x ir=0x%08x opcode=0x%02x rd=%0d rs1=%0d rs2=%0d", dut.cpu_core.pc_ir, dut.cpu_core.ir, dut.cpu_core.opcode, dut.cpu_core.rd, dut.cpu_core.rs1, dut.cpu_core.rs2);
			end

			if (rst_n && dut.wena_mem) begin
				store_count++;
				$display("[STORE] cycle=%0d addr_word=%0d wstrb=0x%0x wdata=0x%08x", cycles, dut.dmem_addr, dut.store_strb, dut.store_wdata);
				if (dut.dmem_addr == stop_addr_word) begin
					last_word0_wdata = dut.store_wdata;
					// PASS: exact match of stop_wdata (default 0xDEADBEEF)
					if (use_stop_wdata && (dut.store_strb == 4'hF) && (dut.store_wdata == stop_wdata)) begin
						saw_store_to_word0 = 1'b1;
					end
					// FAIL: 0xBAD0xxxx (code in low 16 bits)
					else if ((dut.store_strb == 4'hF) && ((dut.store_wdata & 32'hFFFF_0000) == 32'hBAD0_0000)) begin
						saw_store_to_word0 = 1'b1;
						saw_fail_signature = 1'b1;
					end
					// Legacy behavior if someone explicitly disables STOP_WDATA handling.
					else if (!use_stop_wdata && (dut.store_wdata != 32'h0000_0000)) begin
						saw_store_to_word0 = 1'b1;
					end
				end
			end
		end

		if (!saw_store_to_word0) begin
			$fatal(1, "Timeout: no stop store observed within %0d cycles. Default is store 0x%08x to dmem[word %0d]. Optional: +STOP_WDATA=<hex>, +STOP_ADDR=<word>, +MAX_CYCLES=<n>.", max_cycles, stop_wdata, stop_addr_word);
		end
		if (saw_fail_signature) begin
			$fatal(1, "FAIL signature observed at dmem[word %0d]: wdata=0x%08x (code=0x%04x)", stop_addr_word, last_word0_wdata, last_word0_wdata[15:0]);
		end

		// dmem is synchronous; allow the write to commit before reading mem[]
		@(posedge clk);

		$display("---- FINAL SNAPSHOT ----");
		$display("cycles=%0d pc_output=0x%08x cpu_state=%0d ir=0x%08x", cycles, dut.cpu_core.pc_output, dut.cpu_core.cpu_state, dut.cpu_core.ir);
		$display("------------------------");

		dump_dmem();
		$finish;
	end

endmodule

